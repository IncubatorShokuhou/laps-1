netcdf lst {

    dimensions:
        record = unlimited,
        z = 1,
	x = 125,
	y = 105,
        nav = 1,
        namelen = 132;
		
    variables:
        //      lifted index            //

        float
            li(record,z,y,x);
            li:navigation_dim = "nav";
            li:record = "valtime, reftime";
            li:_FillValue = 1.e+37f;
            li:long_name="lifted index";
            li:units="degrees Kelvin";
            li:valid_range= -20000.f, 20000.f;
            li:LAPS_var="LI";
            li:lvl_coord="AGL";
            li:LAPS_units="K";
 
        //      positive buoyant energy         //
        float
            pbe(record,z,y,x);
            pbe:navigation_dim = "nav";
            pbe:record = "valtime, reftime";
            pbe:_FillValue = 1.e+37f;
            pbe:long_name="positive buoyant energy";
            pbe:units="joules/kilogram";
            pbe:valid_range= -20000.f, 20000.f;
            pbe:LAPS_var="PBE";
            pbe:lvl_coord="AGL";
            pbe:LAPS_units="J/KG";
 
         //      negative buoyant energy         //

         float
            nbe(record,z,y,x);
            nbe:navigation_dim = "nav";
            nbe:record = "valtime, reftime";
            nbe:_FillValue = 1.e+37f;
            nbe:long_name="negative buoyant energy";
            nbe:units="joules/kilogram";
            nbe:valid_range= -20000.f, 20000.f;
            nbe:LAPS_var="NBE";
            nbe:lvl_coord="AGL";
            nbe:LAPS_units="J/KG";
 
         //      showalter index        //

         float
            si(record,z,y,x);
            si:navigation_dim = "nav";
            si:record = "valtime, reftime";
            si:_FillValue = 1.e+37f;
            si:long_name="showalter index";
            si:units="degrees kelvin";
            si:valid_range= -20000.f, 20000.f;
            si:LAPS_var="SI";
            si:lvl_coord="AGL";
            si:LAPS_units="K";
 
         //      total totals index         //

         float
            tt(record,z,y,x);
            tt:navigation_dim = "nav";
            tt:record = "valtime, reftime";
            tt:_FillValue = 1.e+37f;
            tt:long_name="total totals index";
            tt:units="degrees kelvin";
            tt:valid_range= -20000.f, 20000.f;
            tt:LAPS_var="TT";
            tt:lvl_coord="AGL";
            tt:LAPS_units="K";
 
         //      k index         //

         float
            k(record,z,y,x);
            k:navigation_dim = "nav";
            k:record = "valtime, reftime";
            k:_FillValue = 1.e+37f;
            k:long_name="k index";
            k:units="degrees kelvin";
            k:valid_range= -20000.f, 20000.f;
            k:LAPS_var="K";
            k:lvl_coord="AGL";
            k:LAPS_units="K";
 
         //      lifted condensation level         //

         float
            lcl(record,z,y,x);
            lcl:navigation_dim = "nav";
            lcl:record = "valtime, reftime";
            lcl:_FillValue = 1.e+37f;
            lcl:long_name="lifted condensation level";
            lcl:units="meters";
            lcl:valid_range= -20000.f, 20000.f;
            lcl:LAPS_var="LCL";
            lcl:lvl_coord="MSL";
            lcl:LAPS_units="M";
 
         //      wet bulb zero         //

         float
            wb0(record,z,y,x);
            wb0:navigation_dim = "nav";
            wb0:record = "valtime, reftime";
            wb0:_FillValue = 1.e+37f;
            wb0:long_name="wet bulb zero";
            wb0:units="meters";
            wb0:valid_range= -20000.f, 20000.f;
            wb0:LAPS_var="WB0";
            wb0:lvl_coord="MSL";
            wb0:LAPS_units="M";
 
         //      wet bulb (1.3C) //

         float
            wb1(record,z,y,x);
            wb1:navigation_dim = "nav";
            wb1:record = "valtime, reftime";
            wb1:_FillValue = 1.e+37f;
            wb1:long_name="wet bulb 1";
            wb1:units="meters";
            wb1:valid_range= -20000.f, 20000.f;
            wb1:LAPS_var="WB1";
            wb1:lvl_coord="MSL";
            wb1:LAPS_units="M";
 
        //	LAPS variables

        long
            imax,
            jmax,
            kmax,
            kdim;

        char
            li_comment(record,z,namelen),
            pbe_comment(record,z,namelen),
            nbe_comment(record,z,namelen),
            si_comment(record,z,namelen),
            tt_comment(record,z,namelen),
            k_comment(record,z,namelen),
            lcl_comment(record,z,namelen),
            wb0_comment(record,z,namelen),
            wb1_comment(record,z,namelen),
            asctime(record,namelen);

			
        //	inventory variables

        short
            li_fcinv(record, z);
            li_fcinv:_FillValue= 0s;
              	
        short
            pbe_fcinv(record, z);
            pbe_fcinv:_FillValue= 0s;
              	
        short
            nbe_fcinv(record, z);
            nbe_fcinv:_FillValue= 0s;
              	
        short
            si_fcinv(record, z);
            si_fcinv:_FillValue= 0s;
              	
        short
            tt_fcinv(record, z);
            tt_fcinv:_FillValue= 0s;
              	
        short
            k_fcinv(record, z);
            k_fcinv:_FillValue= 0s;
              	
        short
            lcl_fcinv(record, z);
            lcl_fcinv:_FillValue= 0s;
              	
        short
            wb0_fcinv(record, z);
            wb0_fcinv:_FillValue= 0s;
              	
        short
            wb1_fcinv(record, z);
            wb1_fcinv:_FillValue= 0s;
              	
        //	list of grid levels

        float 
            level(z);
            level:long_name="level of data";
	    level:units = "hectopascals";
                    	
        //      validtime of the grid 

        double
            valtime(record);
            valtime:long_name = "valid time";
            valtime:units = "seconds since (1970-1-1 00:00:00.0)";

        //      reference time of the process

        double
            reftime(record);
            reftime:long_name = "reference time";
            reftime:units = "seconds since (1970-1-1 00:00:00.0)";

        //      nice name for originating center

        char
            origin_name(namelen);

        //      nice name for process

        char
            process_name(namelen);

        //      nice name for grid description instance
        char
            grid_name(namelen);

        //      basic assumption about earth shape
        char
            earth_shape(namelen);

        // navigation variables using 
        // WMO FM 92-VIII Ext.GRIB specification names
  
        char    grid_type(nav, namelen);
                grid_type:long_name = "GRIB-1 grid type";
  
        char    x_dim(nav, namelen);
                x_dim:long_name = "longitude dimension";
  
        char    y_dim(nav, namelen);
                y_dim:long_name = "latitude dimension";
  
        short   Nx(nav);
                Nx:long_name = "number of x points";
  
        short   Ny(nav);
                Ny:long_name =  "number of y points";
  
        float   La1(nav);
                La1:long_name = "first latitude";
                La1:units = "degrees_north";
  
        float   Lo1(nav);
                Lo1:long_name = "first longitude";
                Lo1:units = "degrees_east" ;
    
        float   LoV(nav);
                LoV:long_name = "orientation of grid" ;
                LoV:units = "degrees_east";
  
        float   Latin1(nav);
                Latin1:long_name = "orientation of grid" ;
                Latin1:units = "degrees_north";

        float   Latin2(nav);
                Latin2:long_name = "orientation of grid" ;
                Latin2:units = "degrees_north";

        float   Dx(nav);
                Dx:long_name = "x grid increment";
                Dx:units = "meters";
  
        float   Dy(nav);
                Dy:long_name = "y grid increment";
                Dy:units = "meters";
  
        // end of navigation variables

        :Conventions = "NUWG";
        :history = "created by LAPS Branch of FSL";
        :record = "valtime, reftime";
        :title = "LAPS lst file - LAPS stability indices ";
        :version = 3;

    data:

        earth_shape     = "spherical radius";
        grid_name       = "LAPS lst file - LAPS stability indices";
        process_name    = "LAPS - Local Analysis and Prediction System";
        x_dim           = "x";
        y_dim           = "y";
}                       
