netcdf liw {

    dimensions:
        record = unlimited,
        z = 1,
	x = 125,
	y = 105,
        nav = 1,
        namelen = 132;
		
    variables:
        //	LAPS Li * 600mb Omega

	float                                  
            liw(record,z,y,x);
            liw:navigation_dim = "nav";
            liw:record = "valtime, reftime";
            liw:_FillValue = 1.e+37f;
            liw:long_name="LAPS li * 600mb omega";
            liw:units="kiloPascals/second";
            liw:valid_range= 0.f, 0.100f;
            liw:LAPS_var="LIW";
            liw:lvl_coord="MSL";
	    liw:LAPS_units="K-PA/S";
                	        
        //	Upslope Component of Moisture Flux

	float                                  
            umf(record,z,y,x);
            umf:navigation_dim = "nav";
            umf:record = "valtime, reftime";
            umf:_FillValue = 1.e+37f;
            umf:long_name="Upslope Component of Moisture Flux";
            umf:units="Meters**2/second";
            umf:valid_range= 0.f, 1000.f;
            umf:LAPS_var="UMF";
            umf:lvl_coord="MSL";
	    umf:LAPS_units="M**2/S";
                	        
        //	LAPS variables

        long
            imax,
            jmax,
            kmax,
            kdim;

        char
            liw_comment(record,z,namelen),
            umf_comment(record,z,namelen),
            asctime(record,namelen);

			
        //	inventory variables

        short
            liw_fcinv(record, z);
            liw_fcinv:_FillValue= 0s;
              	
        short
            umf_fcinv(record, z);
            umf_fcinv:_FillValue= 0s;
              	
        //	list of grid levels

        float 
            level(z);
            level:long_name="level of data";
	    level:units = "hectopascals";
                    	
        //      validtime of the grid 

        double
            valtime(record);
            valtime:long_name = "valid time";
            valtime:units = "seconds since (1970-1-1 00:00:00.0)";

        //      reference time of the process

        double
            reftime(record);
            reftime:long_name = "reference time";
            reftime:units = "seconds since (1970-1-1 00:00:00.0)";

        //      nice name for originating center

        char
            origin_name(namelen);

        //      nice name for process

        char
            process_name(namelen);

        //      nice name for grid description instance
        char
            grid_name(namelen);

        //      basic assumption about earth shape
        char
            earth_shape(namelen);

        // navigation variables using 
        // WMO FM 92-VIII Ext.GRIB specification names
  
        char    grid_type(nav, namelen);
                grid_type:long_name = "GRIB-1 grid type";
  
        char    x_dim(nav, namelen);
                x_dim:long_name = "longitude dimension";
  
        char    y_dim(nav, namelen);
                y_dim:long_name = "latitude dimension";
  
        short   Nx(nav);
                Nx:long_name = "number of x points";
  
        short   Ny(nav);
                Ny:long_name =  "number of y points";
  
        float   La1(nav);
                La1:long_name = "first latitude";
                La1:units = "degrees_north";
  
        float   Lo1(nav);
                Lo1:long_name = "first longitude";
                Lo1:units = "degrees_east" ;
    
        float   LoV(nav);
                LoV:long_name = "orientation of grid" ;
                LoV:units = "degrees_east";
  
        float   Latin1(nav);
                Latin1:long_name = "orientation of grid" ;
                Latin1:units = "degrees_north";

        float   Latin2(nav);
                Latin2:long_name = "orientation of grid" ;
                Latin2:units = "degrees_north";

        float   Dx(nav);
                Dx:long_name = "x grid increment";
                Dx:units = "meters";
  
        float   Dy(nav);
                Dy:long_name = "y grid increment";
                Dy:units = "meters";
  
        // end of navigation variables

        :Conventions = "NUWG";
        :history = "created by LAPS Branch of FSL";
        :record = "valtime, reftime";
        :title = "LAPS liw file - LAPS Li * 600mb Omega";
        :version = 3;

    data:

        earth_shape     = "spherical radius";
        grid_name       = "LAPS liw file - LAPS Li * 600mb Omega";
        process_name    = "LAPS - Local Analysis and Prediction System";
        x_dim           = "x";
        y_dim           = "y";
}                       
