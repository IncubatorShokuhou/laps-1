netcdf narrowband {
dimensions:
	radial = UNLIMITED ; 
	Z_bin = 460 ;
	V_bin = 920 ;
	radarNameLen = 5 ;
	siteNameLen = 132 ;
variables:
	byte Z(radial, Z_bin) ;
		Z:long_name = "Reflectivity" ;
		Z:units = "dBZ" ;
		Z:valid_range = '\2', '\376' ;
		Z:below_threshold = '\0' ;
		Z:range_ambiguous = '\1' ;
		Z:_FillValue = '\377' ;
	byte V(radial, V_bin) ;
		V:long_name = "Velocity" ;
		V:units = "meter/second" ;
		V:valid_range = '\2', '\376' ;
		V:below_threshold = '\0' ;
		V:range_ambiguous = '\1' ;
		V:_FillValue = '\377' ;
	byte W(radial, V_bin) ;
		W:long_name = "Spectrum Width" ;
		W:units = "meter/second" ;
		W:valid_range = '\2', '\376' ;
		W:below_threshold = '\0' ;
		W:range_ambiguous = '\1' ;
		W:_FillValue = '\377' ;
	short elevationNumber ;
		elevationNumber:long_name = "Elevation number" ;
		elevationNumber:units = "count" ;
		elevationNumber:valid_range = 1, 25 ;
	float elevationAngle ;
		elevationAngle:long_name = "Elevation angle" ;
		elevationAngle:units = "degree" ;
		elevationAngle:history = "average of last 20 radialElev" ;
		elevationAngle:valid_range = 0., 90. ;
	short numRadials ;
		numRadials:long_name = "Number of radials" ;
		numRadials:valid_range = 0, 400 ;
	float radialAzim(radial) ;
		radialAzim:long_name = "Radial azimuth angle" ;
		radialAzim:units = "degree" ;
		radialAzim:valid_range = 0., 360. ;
	float radialElev(radial) ;
		radialElev:long_name = "Radial elevation angle" ;
		radialElev:units = "degree" ;
		radialElev:valid_range = 0., 90. ;
	double radialTime(radial) ;
		radialTime:long_name = "Time of radial" ;
		radialTime:units = "seconds since 1970-1-1 00:00:00.00" ;
	char siteName(siteNameLen) ;
		siteName:long_name = "Long name of the radar site" ;
	char radarName(radarNameLen) ;
		radarName:long_name = "Official name of the radar" ;
	float siteLat ;
		siteLat:long_name = "Latitude of site" ;
		siteLat:units = "degrees_north" ;
	float siteLon ;
		siteLon:long_name = "Longitude of site" ;
		siteLon:units = "degrees_east" ;
	float siteAlt ;
		siteAlt:long_name = "Altitude of site above mean sea level" ;
		siteAlt:units = "meter" ;
	short VCP ;
		VCP:long_name = "Volume Coverage Pattern" ;
		VCP:units = "Federal Meteorological Handbook 11 Part A Sec. 4.3" ;
	double esStartTime ;
		esStartTime:long_name = "Start time of elevation scan" ;
		esStartTime:units = "seconds since 1970-1-1 00:00:00.00" ;
	double esEndTime ;
		esEndTime:long_name = "End time of elevation scan" ;
		esEndTime:units = "seconds since 1970-1-1 00:00:00.00" ;
	float unambigRange ;
		unambigRange:long_name = "Unambiguous range" ;
		unambigRange:units = "kilometer" ;
	float firstGateRangeZ ;
		firstGateRangeZ:long_name = "Range to 1st Reflectivity gate" ;
		firstGateRangeZ:units = "kilometer" ;
	float firstGateRangeV ;
		firstGateRangeV:long_name = "Range to 1st Doppler gate" ;
		firstGateRangeV:units = "kilometer" ;
	float gateSizeZ ;
		gateSizeZ:long_name = "Reflectivity gate spacing" ;
		gateSizeZ:units = "kilometer" ;
	float gateSizeV ;
		gateSizeV:long_name = "Doppler gate spacing" ;
		gateSizeV:units = "kilometer" ;
	short numGatesZ ;
		numGatesZ:long_name = "Number of reflectivity gates" ;
		numGatesZ:valid_range = 0, 460 ;
	short numGatesV ;
		numGatesV:long_name = "Number of Doppler gates" ;
		numGatesV:valid_range = 0, 920 ;
	float resolutionV ;
		resolutionV:long_name = "Doppler velocity resolution" ;
		resolutionV:units = "meter/second" ;
	float nyquist ;
		nyquist:long_name = "Nyquist velocity" ;
		nyquist:units = "meter/second" ;
	float calibConst ;
		calibConst:long_name = "System gain calibration constant" ;
		calibConst:units = "dB" ;
		calibConst:valid_range = -50., 50. ;
	float atmosAttenFactor ;
		atmosAttenFactor:long_name = "Atmospheric attenuation factor" ;
		atmosAttenFactor:units = "dB/kilometer" ;
	float powDiffThreshold ;
		powDiffThreshold:long_name = "Range de-aliasing threshold" ;
		powDiffThreshold:units = "dB" ;

// global attributes:
		:history = "Encoded into netCDF by LAPS from narrowband data" ;
		:title = "WSR-88D Narrowband Data" ;
		:Conventions = "NUWG" ;
		:origin = "NOAA/ERL Forecast Systems Laboratory, Boulder, CO" ;
		:version = 1. ;
}
