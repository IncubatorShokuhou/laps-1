netcdf lfr {

    dimensions:
        record = unlimited,
        z = 1,
	x = 125,
	y = 105,
        nav = 1,
        namelen = 132;
		
    variables:
        //	pbl top pressure

	float                                  
            ptp(record,z,y,x);
            ptp:navigation_dim = "nav";
            ptp:record = "valtime, reftime";
            ptp:_FillValue = 1.e+37f;
            ptp:long_name="pbl top pressure";
            ptp:units="pascals";
            ptp:valid_range= 0.f, 10000.f;
            ptp:LAPS_var="PTP";
            ptp:lvl_coord="";
	    ptp:LAPS_units="PA";
                	        
        //	pbl top in meters agl (i.e. depth)
        float 
            pdm(record,z,y,x) ;
            pdm:navigation_dim = "nav";
            pdm:record = "valtime, reftime";
            pdm:_FillValue = 1.e+37f;
            pdm:long_name = "pbl top height" ;
            pdm:units = "meters" ;
            pdm:valid_range = 0.f, 6.0f ;
            pdm:LAPS_var = "PTM" ;
            pdm:lvl_coord = "AGL" ;
            pdm:LAPS_units = "M" ;

        //	LAPS variables

        long
            imax,
            jmax,
            kmax,
            kdim;

        char
            ptp_comment(record,z,namelen),
            pdm_comment(record,z,namelen),
            asctime(record,namelen);

			
        //	inventory variables

        short
            ptp_fcinv(record, z);
            ptp_fcinv:_FillValue= 0s;
              	
        short
            pdm_fcinv(record, z);
            pdm_fcinv:_FillValue= 0s;
              	
        //	list of grid levels

        float 
            level(z);
            level:long_name="level of data";
	    level:units = "hectopascals";
                    	
        //      validtime of the grid 

        double
            valtime(record);
            valtime:long_name = "valid time";
            valtime:units = "seconds since (1970-1-1 00:00:00.0)";

        //      reference time of the process

        double
            reftime(record);
            reftime:long_name = "reference time";
            reftime:units = "seconds since (1970-1-1 00:00:00.0)";

        //      nice name for originating center

        char
            origin_name(namelen);

        //      nice name for process

        char
            process_name(namelen);

        //      nice name for grid description instance
        char
            grid_name(namelen);

        //      basic assumption about earth shape
        char
            earth_shape(namelen);

        // navigation variables using 
        // WMO FM 92-VIII Ext.GRIB specification names
  
        char    grid_type(nav, namelen);
                grid_type:long_name = "GRIB-1 grid type";
  
        char    x_dim(nav, namelen);
                x_dim:long_name = "longitude dimension";
  
        char    y_dim(nav, namelen);
                y_dim:long_name = "latitude dimension";
  
        short   Nx(nav);
                Nx:long_name = "number of x points";
  
        short   Ny(nav);
                Ny:long_name =  "number of y points";
  
        float   La1(nav);
                La1:long_name = "first latitude";
                La1:units = "degrees_north";
  
        float   Lo1(nav);
                Lo1:long_name = "first longitude";
                Lo1:units = "degrees_east" ;
    
        float   LoV(nav);
                LoV:long_name = "orientation of grid" ;
                LoV:units = "degrees_east";
  
        float   Latin1(nav);
                Latin1:long_name = "orientation of grid" ;
                Latin1:units = "degrees_north";

        float   Latin2(nav);
                Latin2:long_name = "orientation of grid" ;
                Latin2:units = "degrees_north";

        float   Dx(nav);
                Dx:long_name = "x grid increment";
                Dx:units = "meters";
  
        float   Dy(nav);
                Dy:long_name = "y grid increment";
                Dy:units = "meters";
  
        // end of navigation variables

        :Conventions = "NUWG";
        :history = "created by LAPS Branch of FSL";
        :record = "valtime, reftime";
        :title = "LAPS pbl file - boundary layer info";
        :version = 3;

    data:

        earth_shape     = "spherical radius";
        grid_name       = "LAPS pbl file - boundary layer info";
        process_name    = "LAPS - Local Analysis and Prediction System";
        x_dim           = "x";
        y_dim           = "y";
}                       
