netcdf lga {

    dimensions:
        record = unlimited,
        z = 21,
	x = 125,
	y = 105,
        nav = 1,
        namelen = 132;
		
    variables:
        //	Background height	

	float                                  
            ht(record,z,y,x);
            ht:navigation_dim = "nav";
            ht:record = "valtime, reftime";
            ht:_FillValue = 1.e+37f;
            ht:long_name="Background height";
            ht:units="meters";
            ht:valid_range= -400.f, 20000.f;
            ht:LAPS_var="HT";
            ht:lvl_coord="SIGMA_P";
	    ht:LAPS_units="METERS";
                	        
        //      Background temperature
 
        float
            t3(record,z,y,x);
            t3:navigation_dim = "nav";
            t3:record = "valtime, reftime";
            t3:_FillValue = 1.e+37f;
            t3:long_name="Background temperature";
            t3:units="degrees Kelvin";
            t3:valid_range= 100.f, 330.f;
            t3:LAPS_var="T3";
            t3:lvl_coord="SIGMA_P";
            t3:LAPS_units="KELVIN";
 

        //      Background specific humidity  //

        float
            sh(record,z,y,x);
            sh:navigation_dim = "nav";
            sh:record = "valtime, reftime";
            sh:_FillValue = 1.e+37f;
            sh:long_name="Background specific humidity";
            sh:units="none";
            sh:valid_range= 0.f, 1.f;
            sh:LAPS_var="SH";
            sh:lvl_coord="SIGMA_P";
            sh:LAPS_units="NONE";
 
        //      Background u wind component   //

        float
            u3(record,z,y,x);
            u3:navigation_dim = "nav";
            u3:record = "valtime, reftime";
            u3:_FillValue= 1.e+37f;
            u3:long_name="Background u wind component";
            u3:units="meters/second";
            u3:valid_range= -200.f, 200.f;
            u3:LAPS_var="U3";
            u3:lvl_coord="SIGMA_P";
            u3:LAPS_units="M/S";
 
        //      Background v wind component           //

        float
            v3(record,z,y,x);
            v3:navigation_dim = "nav";
            v3:record = "valtime, reftime";
            v3:_FillValue= 1.e+37f;
            v3:long_name="Background v wind component";
            v3:valid_range= -200.f, 200.f;
            v3:units="meters/second";
            v3:LAPS_var="V3";
            v3:lvl_coord="SIGMA_P";
            v3:LAPS_units="M/S";
 
        //      Background w wind component           //

        float
            om(record,z,y,x);
            om:navigation_dim = "nav";
            om:record = "valtime, reftime";
            om:_FillValue= 1.e+37f;
            om:long_name="Background w wind component";
            om:valid_range= -100.f, 100.f;
            om:units="pascals/second";
            om:LAPS_var="OM";
            om:lvl_coord="SIGMA_P";
            om:LAPS_units="PA/S";
 

        //	LAPS variables

        long
            imax,
            jmax,
            kmax,
            kdim;

        char
            ht_comment(record,z,namelen),
            t3_comment(record,z,namelen),
            sh_comment(record,z,namelen),
            u3_comment(record,z,namelen),
            v3_comment(record,z,namelen),
            om_comment(record,z,namelen),
            asctime(record,namelen);

			
        //	inventory variables

        short
            ht_fcinv(record, z);
            ht_fcinv:_FillValue= 0s;
              	
        short
            t3_fcinv(record, z);
            t3_fcinv:_FillValue= 0s;
              	
        short
            sh_fcinv(record, z);
            sh_fcinv:_FillValue= 0s;
              	
        short
            u3_fcinv(record, z);
            u3_fcinv:_FillValue= 0s;
              	
        short
            v3_fcinv(record, z);
            v3_fcinv:_FillValue= 0s;
              	
        short
            om_fcinv(record, z);
            om_fcinv:_FillValue= 0s;
              	
        //	list of grid levels

        float 
            level(z);
            level:long_name="level of data";
	    level:units = "hectopascals";
                    	
        //      validtime of the grid 

        double
            valtime(record);
            valtime:long_name = "valid time";
            valtime:units = "seconds since (1970-1-1 00:00:00.0)";

        //      reference time of the process

        double
            reftime(record);
            reftime:long_name = "reference time";
            reftime:units = "seconds since (1970-1-1 00:00:00.0)";

        //      nice name for originating center

        char
            origin_name(namelen);

        //      nice name for process

        char
            process_name(namelen);

        //      nice name for grid description instance
        char
            grid_name(namelen);

        //      basic assumption about earth shape
        char
            earth_shape(namelen);

        // navigation variables using 
        // WMO FM 92-VIII Ext.GRIB specification names
  
        char    grid_type(nav, namelen);
                grid_type:long_name = "GRIB-1 grid type";
  
        char    x_dim(nav, namelen);
                x_dim:long_name = "longitude dimension";
  
        char    y_dim(nav, namelen);
                y_dim:long_name = "latitude dimension";
  
        short   Nx(nav);
                Nx:long_name = "number of x points";
  
        short   Ny(nav);
                Ny:long_name =  "number of y points";
  
        float   La1(nav);
                La1:long_name = "first latitude";
                La1:units = "degrees_north";
  
        float   Lo1(nav);
                Lo1:long_name = "first longitude";
                Lo1:units = "degrees_east" ;
    
        float   LoV(nav);
                LoV:long_name = "orientation of grid" ;
                LoV:units = "degrees_east";
  
        float   Latin1(nav);
                Latin1:long_name = "orientation of grid" ;
                Latin1:units = "degrees_north";

        float   Latin2(nav);
                Latin2:long_name = "orientation of grid" ;
                Latin2:units = "degrees_north";

        float   Dx(nav);
                Dx:long_name = "x grid increment";
                Dx:units = "meters";
  
        float   Dy(nav);
                Dy:long_name = "y grid increment";
                Dy:units = "meters";
  
        // end of navigation variables

        :Conventions = "NUWG";
        :history = "created by LAPS Branch of FSL";
        :record = "valtime, reftime";
        :title = "LAPS lga file - background analysis fields";
        :version = 3;

    data:

        earth_shape     = "spherical radius";
        grid_name       = "LAPS lga file - background analysis fields";
        process_name    = "LAPS - Local Analysis and Prediction System";
        x_dim           = "x";
        y_dim           = "y";
}                       
